`timescale 1ns/1ns

// Creacion del modulo
module MEM
(
	input MEM_WRITE, // WRITE / READ
	input [31:0]WRITE_DATA, // Dato
	output reg [31:0]READ_DATA, // Salida (Si estamos leyendo)
	input [31:0]ADRESS // Direccion donde estamos apuntando
);

// Registro / Cables
reg [31:0] memory [31:0]; // <-- Memoria

// Bloque always
always @*
begin
	if (MEM_WRITE) // Si es modo WRITE
	begin
		memory[ADRESS] = WRITE_DATA; // <-- Escribir
		READ_DATA = 32'dx;
	end
	else // Si no, es modo READ
	begin
		READ_DATA = memory[ADRESS]; // <-- Leer
	end
end

endmodule : MEM